library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
USE work.aux_package.all;
---------------------------------------------------------
entity tb_datapath is
	constant n : integer := 8;
end tb_datapath;
---------------------------------------------------------
architecture rtb of tb_datapath is
	signal clk,rst,ena : std_logic;
signal	mov, st,ld, jnc, jc ,jmp, sub, add,nop, Nflag, Zflag,Cflag,Cout, Cin, Ain, RFin, RFout,IRin,PCin,Imm1_in,Imm2_in,done_in,DoneProgram,Mem_wr, Mem_out, Mem_in		 : std_logic;
signal	OPC															: std_logic_vector(3 downto 0);
signal	RFadder ,PCsel												: std_logic_vector(1 downto 0);
signal  DataMemTBDataIn,ProgMemTBDataIn	,DataMemDataOut 			: std_logic_vector(16-1 downto 0);
signal	ProgMemTBWren				 	 							:  std_logic;
signal	DataMemTBWren 												:  std_logic;
signal	ProgMemTbWAddr												: std_logic_vector(6-1 downto 0);
signal	DataMemTbWAddr,DataMemTbRAddr								: std_logic_vector(6-1 downto 0);
signal	TBactive           											: std_logic;
	
	
begin
	DataPath1		: Datapath 	generic map (16, 6,4, 64)   port map(rst,clk,mov,st,ld,done_in,  jnc, jc ,jmp, sub, add,nop, Nflag, Zflag,Cflag
																			  ,Cout, Cin, Ain, RFin, RFout,IRin,PCin,Imm1_in,Imm2_in,Mem_wr, Mem_out, Mem_in,
																			  OPC,RFadder ,PCsel,ProgMemTBDataIn,DataMemTBDataIn,DataMemDataOut,ProgMemTBWren=>ProgMemTBWren,DataMemTBWren=>DataMemTBWren,ProgMemTbWAddr=>ProgMemTbWAddr,DataMemTbRAddr=>DataMemTbRAddr,DataMemTbWAddr=>DataMemTbWAddr,TBactive=>TBactive);

	--------- start of stimulus section ------------------	
	DataMemTbRAddr <= (others => '0');
        gen_clk : process
        begin
		  clk <= '0';
		  wait for 50 ns;
		  clk <= not clk;
		  wait for 50 ns;
        end process;
		gen_memorey : process
		variable    TempWAddresses		: std_logic_vector(5 downto 0) ;
		variable    TempWData			: std_logic_vector(15 downto 0) ;
		variable    TempWprog			: std_logic_vector(15 downto 0) ;
		variable 	counter				: integer;

        begin
		  TempWAddresses := (others => '0');
		  TempWData      :=	(others => '0');		
		  counter := 0;	 
		  rst <='1';
		  TBactive <= '0';
		  DataMemTBWren <= '1';
		  ProgMemTBWren <= '1';
		while counter < 15 loop
			if counter = 0 then 
				TempWprog      :=	"1001000100000001";			--ld
			elsif counter = 1 then  
				TempWprog      := 	"1001001000000111";			--ld
			elsif counter = 2 then  
				TempWprog      := 	"0000011000010010";--add r6 <- r2+r1
			elsif counter = 3 then  
				TempWprog      := 	"0001000101100010";	--sub r1 = r6-r2
			elsif counter = 4 then  
				TempWprog      := 	"0010110000110010";		--nop
			elsif counter = 5 then  
				TempWprog      := 	"0100000000000000";	-- jmp offset 0
			elsif counter = 6 then  
				TempWprog      := 	"0101000000000001";		-- jc 1
			elsif counter = 7 then  
				TempWprog      := 	"0110000000000011"; -- jnc 3
			elsif counter = 8 then  
				TempWprog      := 	"1000111100110010"; --mov r15 <- 00110010
			elsif counter = 9 then  
				TempWprog      := 	"0001000100010010";		-- sub r1 = r1-r2		
			elsif counter = 10 then  
				TempWprog      := 	"0100111111111101";			 -- jmp -3		
			elsif counter = 11 then  
				TempWprog      := 	"1010000100001100"; -- str [r0+12] <- r1
			elsif counter = 12 then  
				TempWprog      := 	"1010001000111100";	-- str [r3+12] <- r2
			elsif counter = 13 then  
				TempWprog      := 	"1010111100101101"; -- str [r2+13] <- r15
			elsif counter = 14 then  
				TempWprog      := 	"1010011001101111";-- str [r6+15] <- r6
			end if;
			DataMemTbWAddr <= TempWAddresses;
			ProgMemTbWAddr <= TempWAddresses;
			ProgMemTBDataIn <= TempWprog ;
			DataMemTBDataIn <= TempWData;
			wait until rising_edge(clk);
			TempWAddresses := TempWAddresses +1;
			TempWData      :=	TempWData + 1;
			counter := counter + 1;
		end loop ;
			rst <='0';
			TBactive <= '1';
			DataMemTBWren <= '0';
			ProgMemTBWren <= '0';
		wait;
        end process;
	
		gen_input : process
		variable 	counter			: integer;
        begin
		counter := 0;
		wait until rst = '0' and TBactive = '1';
		
		while counter < 71 loop 
			ena <= '1';
			if counter = 0  then --fecth ld1 
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 1  then -- decode ld1
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 2  then --cyc 1 ld 1
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 3  then --cyc 2 ld1
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='1';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 4  then -- cyc 3 ld1
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '1';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";
			elsif counter = 5  then -- cyc 4 ld1
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0'; 
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';  
				Mem_out <= '1'; 
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";	
			elsif counter = 6  then --fecth ld2
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 7  then --decode ld2
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 8  then --cyc 1 ld2
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 9  then --cyc 2 ld2
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='1';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 10  then --cyc 3 ld2
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '1';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";
			elsif counter = 11  then --cyc 4 ld2
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0' ;
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0'  ;
				Mem_out <= '1' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
			elsif counter = 12  then  --fecth add 
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 13  then --decode add
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 14  then --cyc 1 add
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 15  then--cyc 2 add
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 16  then --cyc 3 add
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
			elsif counter = 17  then--fecth sub
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0' ;
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0' ; 
				Mem_out <= '0' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
			elsif counter = 18  then --decode sub
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 19  then --cyc 1 sub
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";	
							
			elsif counter = 20  then--cyc 2 sub
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0001";
				RFadder<="00";
				PCsel  <="00";														
				
			elsif counter = 21  then--cyc 3 sub
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0001";
				RFadder<="10";
				PCsel  <="10";

			elsif counter = 22  then--fecth nop
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0' ;
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0' ; 
				Mem_out <= '0' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
			elsif counter = 23  then--decode nop
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 24  then--cyc1 nop
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";	
							
			elsif counter = 25  then--cyc2 nop
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0001";
				RFadder<="00";
				PCsel  <="00";														
				
			elsif counter = 26  then--cyc3 nop
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0001";
				RFadder<="10";
				PCsel  <="10";				
			elsif counter = 27 then -- fecth jmp 0
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 28  then -- decode jmp 0
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 29  then --excute jmp 0
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='1';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="01";	
			elsif counter = 30 then-- fecth jc 1
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
				
			elsif counter = 31  then-- fecth jc 1
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";		
				
			elsif counter = 32  then-- excute jc 1
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='1';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				if Cflag = '1' then
					PCsel  <="01";
				else
					PCsel  <="10";
				end if;
			elsif counter = 33 then -- fecth mov 
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
				
			elsif counter = 34  then -- decode mov 
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";		
				
			elsif counter = 35  then --excute mov r15 <- 00110010
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0' ;
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='1';
				Imm2_in <='0';
				Mem_wr <= '0'  ;
				Mem_out <= '0' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
				
			elsif counter = 36  then  --fecth sub
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 37  then --decode sub
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 38  then --cyc 1 sub
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 39  then--cyc 2 sub
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0001";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 40  then --cyc 3 sub
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='1';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
			elsif counter = 41 then -- fecth jmp -3
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 42  then -- decode jmp -3
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 43  then --excute jmp -3
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='1';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="01";					
			elsif counter = 44 then-- fecth jnc 3
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
				
			elsif counter = 45  then-- decode jnc 3
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";		
				
			elsif counter = 46  then-- excute jnc 3
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='1';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				if Cflag = '0' then
					PCsel  <="01";
				else
					PCsel  <="10";
				end if;
			elsif counter = 47  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 48  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 49  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 50  then
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='1';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 51  then
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '1';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";
			elsif counter = 52  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1' ;
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '1'  ;
				Mem_out <= '0' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
			elsif counter = 53  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 54  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 55  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 56  then
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='1';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 57  then
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '1';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";
			elsif counter = 58  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1' ;
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '1'  ;
				Mem_out <= '0' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
			elsif counter = 59  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 60  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 61  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 62  then
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='1';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 63  then
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '1';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";
			elsif counter = 64  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1' ;
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '1'  ;
				Mem_out <= '0' ;
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";
			elsif counter = 65  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';
				RFin   <='0';
				RFout  <='0';
				IRin   <='1';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";
			elsif counter = 66  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 67  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '1';						
				RFin   <='0';
				RFout  <='1';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
    			Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";														
				
			elsif counter = 68  then
				cout 	<= '0';
				cin		<= '1';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='1';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="00";
				PCsel  <="00";	
							
			elsif counter = 69  then
				cout 	<= '1';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='0';
				IRin   <='0';
				PCin   <='0';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '0';
				Mem_out <= '0';
				Mem_in <= '1';
				OPC    <="0000";
				RFadder<="01";
				PCsel  <="00";
			elsif counter = 70  then
				cout 	<= '0';
				cin		<= '0';
				Ain		<= '0';						
				RFin   <='0';
				RFout  <='1'; 
				IRin   <='0';
				PCin   <='1';
				Imm1_in <='0';
				Imm2_in <='0';
				Mem_wr <= '1' ; 
				Mem_out <= '0'; 
				Mem_in <= '0';
				OPC    <="0000";
				RFadder<="10";
				PCsel  <="10";				
	

			end if;
			wait until rising_edge(clk);
			counter := counter + 1;
		end loop ;
		ena <= '0';
		wait;
        end process;		

		
				
end architecture rtb;
